/***********************************************************************/
/*********            		 	XXXX.sv     	    	 	************/
/*********                   V1.0(20160000)					************/
/*********           Written By Morning---20160718          ************/
/***********************************************************************/


/*=====================================================================*/

/*----------------------------block function---------------------------*/

/*=====================================================================*/






/*---------------------------------------------------------------------*/



/*=====================================================================*/



//=======================================================================
//--------------------------End of XXXXXXXX.sv---------------------------
//=======================================================================
